module Core(
  input   clock,
  input   reset
);
endmodule
